module myModule();

initial
 begin
  $display("hello world");
  $finish;
 end
endmodule

